module negate(in, out);
  input in
  output out
  assign out != in //unsure if correct?
    
    endmodule :negate;
