`timescale 1ns / 1ps

module logicalNot(output [31:0]out, input [31:0]in);

  assign out = ~in; 
    
endmodule 
