`timescale 1ns / 1ps

module logicalAnd(input [31:0] in2, in1, output [31:0]out);

assign out = in1 & in2;

endmodule
