`timescale 1ns / 1ps

module logicalNot(output out[31:0], input in[31:0]);

  assign out = ~in; 
    
endmodule 
